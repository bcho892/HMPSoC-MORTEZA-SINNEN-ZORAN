-- zoran_nios_biglari_sseg_0.vhd

-- Generated using ACDS version 18.1 646

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity zoran_nios_biglari_sseg_0 is
	port (
		done          : out std_logic;                                        -- nios_custom_instruction_slave.done
		clock         : in  std_logic                     := '0';             --                              .clk
		display_value : in  std_logic_vector(31 downto 0) := (others => '0'); --                              .dataa
		start         : in  std_logic                     := '0';             --                              .start
		hex0          : out std_logic_vector(6 downto 0);                     --                   conduit_end.zoran0
		hex1          : out std_logic_vector(6 downto 0);                     --                              .zoran1
		hex2          : out std_logic_vector(6 downto 0);                     --                              .zoran2
		hex3          : out std_logic_vector(6 downto 0);                     --                              .zoran3
		hex4          : out std_logic_vector(6 downto 0);                     --                              .zoran4
		hex5          : out std_logic_vector(6 downto 0)                      --                              .zoran5
	);
end entity zoran_nios_biglari_sseg_0;

architecture rtl of zoran_nios_biglari_sseg_0 is
	component ci_read_item_instruction is
		port (
			done          : out std_logic;                                        -- done
			clock         : in  std_logic                     := 'X';             -- clk
			display_value : in  std_logic_vector(31 downto 0) := (others => 'X'); -- dataa
			start         : in  std_logic                     := 'X';             -- start
			hex0          : out std_logic_vector(6 downto 0);                     -- zoran0
			hex1          : out std_logic_vector(6 downto 0);                     -- zoran1
			hex2          : out std_logic_vector(6 downto 0);                     -- zoran2
			hex3          : out std_logic_vector(6 downto 0);                     -- zoran3
			hex4          : out std_logic_vector(6 downto 0);                     -- zoran4
			hex5          : out std_logic_vector(6 downto 0)                      -- zoran5
		);
	end component ci_read_item_instruction;

begin

	biglari_sseg_0 : component ci_read_item_instruction
		port map (
			done          => done,          -- nios_custom_instruction_slave.done
			clock         => clock,         --                              .clk
			display_value => display_value, --                              .dataa
			start         => start,         --                              .start
			hex0          => hex0,          --                   conduit_end.zoran0
			hex1          => hex1,          --                              .zoran1
			hex2          => hex2,          --                              .zoran2
			hex3          => hex3,          --                              .zoran3
			hex4          => hex4,          --                              .zoran4
			hex5          => hex5           --                              .zoran5
		);

end architecture rtl; -- of zoran_nios_biglari_sseg_0
