-- This file should be updated using the script called generate_file_paths.py at the root
package FilePaths is
   constant RECOP_FIXED_CONFIG_FILE_PATH : string := "C:\Users\AKLbc\Desktop\Development\HMPSoC-MORTEZA-SINNEN-ZORAN\src\recop_programs\configuration.mif";
   constant RECOP_CONFIGURABLE_CONFIG_FILE_PATH : string := "C:\Users\AKLbc\Desktop\Development\HMPSoC-MORTEZA-SINNEN-ZORAN\src\recop_programs\user_configuration.mif";
   constant RECOP_VALUED_CONFIG_FIELDS_FILE_PATH : string := "C:\Users\AKLbc\Desktop\Development\HMPSoC-MORTEZA-SINNEN-ZORAN\src\recop_programs\valued_config_fields.mif";
   constant RECOP_WOLF_CONFIG_FIELDS_FILE_PATH : string := "C:\Users\AKLbc\Desktop\Development\HMPSoC-MORTEZA-SINNEN-ZORAN\src\recop_programs\config_core_window.mif";
end package;