library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;

package FilePaths is
    constant RECOP_FIXED_CONFIG_FILE_PATH         : string := "C:\Users\AKLbc\Desktop\Development\HMPSoC-MORTEZA-SINNEN-ZORAN\src\recop_programs\configuration.mif";
    constant RECOP_CONFIGURABLE_CONFIG_FILE_PATH  : string := "C:\Users\AKLbc\Desktop\Development\HMPSoC-MORTEZA-SINNEN-ZORAN\src\recop_programs\user_configuration.mif";
    constant RECOP_VALUED_CONFIG_FIELDS_FILE_PATH : string := "H:\Documents\GitHub\701-hmpsoc\HMPSoC-MORTEZA-SINNEN-ZORAN\src\recop_programs\valued_config_fields";
end package;