library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;

package FilePaths is
    constant RECOP_FILE_PATH : string := "C:\Users\AKLbc\Desktop\Development\HMPSoC-MORTEZA-SINNEN-ZORAN\src\recop_programs\configuration.mif";
end package;